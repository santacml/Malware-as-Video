module DE1_SoC (
	    CLOCK_50,
	    KEY,
	    SW,
	    HEX0,
	    HEX1,
	    HEX2,
	    HEX3,
	    HEX4,
	    HEX5,
	    LEDR,
		UART_RXD,
		UART_TXD

	    );

   input CLOCK_50;
   input [3:0] KEY;
   input [9:0] SW;
   output [6:0] HEX0, HEX1,  HEX2,  HEX3,  HEX4,  HEX5;
   reg [6:0] 	hex0, hex1, hex2, hex3, hex4, hex5, hex6, hex7;
   
   integer clkCount = 0;
   reg clkDone = 0;
   
   output [7:0] LEDR;
    input UART_RXD;
    output UART_TXD;    
	wire clk = CLOCK_50;
	wire go = ~KEY[1];


   wire 	reset = ~KEY[0];
   wire 	start;
   wire [31:0] 	return_val;
   reg  [31:0] 	return_val_reg;
   wire 	finish;
   wire [3:0]	state;

   //hex_digits h7( .x(hex7), .hex_LEDs(HEX7));
   //hex_digits h6( .x(hex6), .hex_LEDs(HEX6));
   hex_digits h5( .x(hex5), .hex_LEDs(HEX5));
   hex_digits h4( .x(hex4), .hex_LEDs(HEX4));
   hex_digits h3( .x(hex3), .hex_LEDs(HEX3));
   hex_digits h2( .x(hex2), .hex_LEDs(HEX2));
   hex_digits h1( .x(hex1), .hex_LEDs(HEX1));
   hex_digits h0( .x(hex0), .hex_LEDs(HEX0));
   
	always @ (*) begin
		hex5 <= return_val_reg;
		hex4 <= y_Q;
                hex3 <= clk;
	end
    assign UART_TXD = 1'b0;

    parameter s_WAIT = 3'b001, s_START = 3'b010, s_EXE = 3'b011,
                s_DONE = 3'b100;

    // state registers
    reg [3:0] y_Q, Y_D;

    assign LEDR[3:0] = y_Q;

    // next state
    always @(*)
    begin
        case (y_Q)
            s_WAIT: if (go) Y_D = s_START; else Y_D = y_Q;

            s_START: Y_D = s_EXE;

            s_EXE: if (!finish) Y_D = s_EXE; else Y_D = s_DONE;

            s_DONE: Y_D = s_DONE;

            default: Y_D = 3'bxxx;
        endcase
    end

    // current state
    always @(posedge clk)
    begin

	if (reset) begin // synchronous clear
            y_Q <= s_WAIT;
	    hex2 <= 0;
	    hex1 <= 0;
	    hex0 <= 0;
	end
        else
            y_Q <= Y_D;

    end
	
    always @(posedge clk)
	if (y_Q == s_EXE && (!finish))
            clkCount <= clkCount + 1;
        else if (y_Q == s_EXE && finish && (0 == clkDone)) begin
            return_val_reg <= return_val;
            clkDone <= 1;
	    //hex3 <= clkCount / 150000000; //seconds (this will be 0, doesn't matter)
            hex2 <= clkCount / 5000000;  //hundreds of ms (casts to int)
            hex1 <=  ((clkCount - clkCount / 5000000) / 500000);   //tens of ms (casts to int)
            hex0 <= ((clkCount - clkCount / 5000000 -  clkCount/ 500000) / 50000);    //single digits ms (casts to int)
         end
        else if (y_Q == s_EXE && finish)
            return_val_reg <= return_val;
        else if (y_Q == s_DONE)
            return_val_reg <= return_val_reg;
        else
            return_val_reg <= 0;



    assign start = (y_Q == s_START);

   
   top top_inst (
      .clk (clk),
      .reset (reset),
      .finish (finish),
      .return_val (return_val),
        .start (start)

    );

endmodule
